* a simple RLC line ckt
Vin 1 0 PWL 0 5.0e-10 2.0 2e-9 2.0 2.5e-9 0 
R_1 1 2 10
L_1 2 3 2e-010
C_1 3 0 1e-013
R_2 3 4 10
L_2 4 5 2e-010
C_2 5 0 1e-013
R_3 5 6 10
L_3 6 7 2e-010
C_3 7 0 1e-013
R_4 7 8 10
L_4 8 9 2e-010
C_4 9 0 1e-013
R_5 9 10 10
L_5 10 11 2e-010
C_5 11 0 1e-013
R_6 11 12 10
L_6 12 13 2e-010
C_6 13 0 1e-013
R_7 13 14 10
L_7 14 15 2e-010
C_7 15 0 1e-013
R_8 15 16 10
L_8 16 17 2e-010
C_8 17 0 1e-013
R_9 17 18 10
L_9 18 19 2e-010
C_9 19 0 1e-013
R_10 19 20 10
L_10 20 21 2e-010
C_10 21 0 1e-013
R_11 21 22 10
L_11 22 23 2e-010
C_11 23 0 1e-013
R_12 23 24 10
L_12 24 25 2e-010
C_12 25 0 1e-013
R_13 25 26 10
L_13 26 27 2e-010
C_13 27 0 1e-013
R_14 27 28 10
L_14 28 29 2e-010
C_14 29 0 1e-013
R_15 29 30 10
L_15 30 31 2e-010
C_15 31 0 1e-013
R_16 31 32 10
L_16 32 33 2e-010
C_16 33 0 1e-013
R_17 33 34 10
L_17 34 35 2e-010
C_17 35 0 1e-013
R_18 35 36 10
L_18 36 37 2e-010
C_18 37 0 1e-013
R_19 37 38 10
L_19 38 39 2e-010
C_19 39 0 1e-013
.TRAN TR 1.0e-11 3e-9
.PLOTNV 2
.PLOTNV 10
.PLOTNV 20
.PLOTNV 39
.end 
