* transmission gate mux

VDD 103 0 DC 3
Vin 101 0 PWL 0 5.0e-10 3.0 0.5e-8 3.0 0.6e-8 0.0 1e-8 0.0 1.1e-8 3.0
Rin 101 102 10
M1 108 102 103 p 30e-6 0.35e-6 1
M2 108 102 0 n 10e-6 0.35e-6 2
Va 100 0 DC 3
Vb 99 0 DC 0

Map 100 102 104 p 60e-6 0.35e-6 1 
Man 100 108 104 n 20e-6 0.35e-6 2 
Mbp 99 108 104 p 60e-6 0.35e-6 1 
Mbn 99 102 104 n 20e-6 0.35e-6 2 

M3 107 104 103 p 30e-6 0.35e-6 1
M4 107 104 0 n 10e-6 0.35e-6 2
C1 107 0 0.1e-12
.MODEL 1 VT -0.75 MU 5e-2 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.MODEL 2 VT 0.83 MU 1.5e-1 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.TRAN TR 1.0e-11 2.0e-8
.PLOTNV 102
.PLOTNV 108
.PLOTNV 104
.PLOTNV 107

