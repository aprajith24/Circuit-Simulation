* simple clock tree contains one driver and three leaf nodes

VDD 103 0 DC 3
Vin 101 0 PWL 0 5.0e-10 3.0
Rin 101 102 10
M11 104 102 103 p 90e-6 0.35e-6 1
M21 104 102 0 n 30e-6 0.35e-6 2
C11 104 0 0.1e-12
R21 104 105 25 
L11 105 106 0.1e-9
C21 106 0 0.9e-12
R22 106 107 25 
L12 107 108 0.1e-9
C22 108 0 0.1e-12
R23 106 109 25 
L13 109 110 0.1e-9
C23 110 0 0.1e-12
R24 106 111 150
L14 111 112 0.6e-9
C24 112 0 0.6e-12
M12 113 108 103 p 60e-6 0.35e-6 1
M22 113 108 0 n 20e-6 0.35e-6 2
M13 114 110 103 p 30e-6 0.35e-6 1
M23 114 110 0 n 10e-6 0.35e-6 2
M14 115 112 103 p 30e-6 0.35e-6 1
M24 115 112 0 n 10e-6 0.35e-6 2
C91 113 0 0.5e-12
C92 114 0 0.5e-12
C93 115 0 0.5e-12
.MODEL 1 VT -0.75 MU 5e-2 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.MODEL 2 VT 0.83 MU 1.5e-1 COX 0.3e-4 LAMBDA 0.05 CJ0 4.0e-14
.TRAN TR 1.0e-11 2.0e-8
.PLOTNV 104
.PLOTNV 106
.PLOTNV 108
.PLOTNV 110
.PLOTNV 112
.PLOTNV 113
.PLOTNV 114
.PLOTNV 115
